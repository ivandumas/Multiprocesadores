module sumador(
    input logic [8:0] absoluto,
    input logic [31:0] sumreg_out,
    output logic [31:0] result
);

assign result = absoluto + sum_out;

endmodule