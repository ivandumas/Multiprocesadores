module controlunit (
    ports
);
    
endmodule