module alu  (
	input  logic [15:0]	A,
	input  logic [15:0]	B,
	input  logic			s0,
	output logic [15:0]	OUT
	);
		
	
	always_comb OUT = s0 ? A + B :  A - B;
					
endmodule
