module ALUcontrol (
    input logic [5:0] func,
    input logic [1:0] ALUOp,
    output logic [2:0] ALUCtrl
);
    
endmodule