module mips (
    
);

endmodule